package test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    import my_env_pkg::*;

    `include "base_test.sv"
endpackage
interface reset_if(
        input  logic clk,
        output logic reset
    );

endinterface